// File: variables.vh
// VARIABLES for IMEM AND DMEM

`ifndef VARIABLES
`define VARIABLES

`define MEM_BYTES_DMEM 64
`define MEM_BYTES_IMEM 256

`endif