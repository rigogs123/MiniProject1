//This module concatenates immediates based on the instruction type and the operation

module imm_gen (
    input wire [4:0] a,
    input wire [4:0] b,
    input wire [10:0] c,
    input wire [1:0] imm_sel_in,
    output wire [31:0] out
);
    


endmodule
