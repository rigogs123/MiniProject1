// File: variables.vh
// VARIABLES for IMEM AND DMEM

`ifndef OPCODES
`define OPCODES

`define R_TYPE 2'b00
`define I_TYPE 2'b01
`define M_TYPE 2'b01
`define B_TYPE 2'b11

`define ADD 4'b0000
`define SUB 4'b0001

`endif