// File: variables.vh
// VARIABLES for IMEM AND DMEM

`ifndef VARIABLES
`define VARIABLES

`define MEM_BYTES_DMEM 32
`define MEM_BYTES_IMEM 32

`endif